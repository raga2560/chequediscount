<div class="panel panel-primary">
                        <div class="panel-heading">
                            Market
							<button  class="btn btn-default" ng-click="refreshmarket()">Refresh Market</button>
                        </div>
                        <div class="panel-body">
<table ng-table="tableParams" class="table" show-filter="true">
    <tr ng-repeat="record in $data">
        <td title="'Issuer'" filter="{ name: 'text'}" sortable="'issuer'">
            {{record.issuer}}</td>
        <td title="'Amount'" filter="{ amount: 'number'}" sortable="'amount'">
            {{record.amount}}</td>
		<td title="'Rating/NW Rating'" filter="{ issuerrating: 'number'}" sortable="'issuerrating'">
		<button class="btn btn-info btn-lg" ng-show="record.issuerrating" >{{record.issuerrating}} /{{record.networkrating}} </button>
            </td>
		<td title="'Discount'" filter="{ discount: 'number'}" sortable="'discount'">
		<button class="btn btn-info btn-lg" ng-show="record.discount" >{{record.discount}} % </button>
            </td>
		<td title="'Exposure'" filter="{ exposure: 'number'}" sortable="'exposure'" ng-show="record.exposure">
            {{record.exposure}} %</td>
		<td title="'IssuerLimit'" filter="{ issuerlimit: 'number'}" sortable="'issuerlimit'">
            {{record.issuerlimit}}</td>
		<td title="'Discounter'" filter="{ discounter: 'text'}" sortable="'discounter'">
            {{record.discounter}}</td>
    </tr>
</table>

</div>
</div>
